//commit 16ae9ddcda54fc9a2fddffad73174cf793ac7814
//Author: Tang Haojin <tanghaojin@outlook.com>
//Date:   Thu Apr 3 22:44:20 2025 +0800
//
//    feat(Top): make address spaces of seperate TL port configurable (#4496)
//    
//    - `SeperateTLBus` and `SeperateTLBusRanges`: Generate a separate
//      TileLink bus with corresponding address ranges
//      - with `XSNoCTopConfig`: Multiple ranges can be specified, and
//        `SeperateDM` is ignored
//      - without `XSNoCTopConfig`: exactly one address range can be specified,
//        and can only be used to connected with DM by `SeperateDM`
//diff --git a/difftest b/difftest
//--- a/difftest
//+++ b/difftest
//@@ -1 +1 @@
//-Subproject commit 62e4540c03c03aa947bdb67f4b6bf66f1a29c5d0
//+Subproject commit 62e4540c03c03aa947bdb67f4b6bf66f1a29c5d0-dirty
// Generated by CIRCT firtool-1.62.1
// Standard header to adapt well known macros for register randomization.
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_MEM_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_MEM_INIT
`endif // not def RANDOMIZE
`ifndef RANDOMIZE
  `ifdef RANDOMIZE_REG_INIT
    `define RANDOMIZE
  `endif // RANDOMIZE_REG_INIT
`endif // not def RANDOMIZE

// RANDOM may be set to an expression that produces a 32-bit random unsigned value.
`ifndef RANDOM
  `define RANDOM $random
`endif // not def RANDOM

// Users can define INIT_RANDOM as general code that gets injected into the
// initializer block for modules with registers.
`ifndef INIT_RANDOM
  `define INIT_RANDOM
`endif // not def INIT_RANDOM

// If using random initialization, you can also define RANDOMIZE_DELAY to
// customize the delay used, otherwise 0.002 is used.
`ifndef RANDOMIZE_DELAY
  `define RANDOMIZE_DELAY 0.002
`endif // not def RANDOMIZE_DELAY

// Define INIT_RANDOM_PROLOG_ for use in our modules below.
`ifndef INIT_RANDOM_PROLOG_
  `ifdef RANDOMIZE
    `ifdef VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM
    `else  // VERILATOR
      `define INIT_RANDOM_PROLOG_ `INIT_RANDOM #`RANDOMIZE_DELAY begin end
    `endif // VERILATOR
  `else  // RANDOMIZE
    `define INIT_RANDOM_PROLOG_
  `endif // RANDOMIZE
`endif // not def INIT_RANDOM_PROLOG_

// Include register initializers in init blocks unless synthesis is set
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_REG_
    `define ENABLE_INITIAL_REG_
  `endif // not def ENABLE_INITIAL_REG_
`endif // not def SYNTHESIS

// Include rmemory initializers in init blocks unless synthesis is set
`ifndef SYNTHESIS
  `ifndef ENABLE_INITIAL_MEM_
    `define ENABLE_INITIAL_MEM_
  `endif // not def ENABLE_INITIAL_MEM_
`endif // not def SYNTHESIS

module SimTop(
  input         clock,
  input         reset,
  output [63:0] difftest_exit,
  output [63:0] difftest_step,
  input         difftest_perfCtrl_clean,
  input         difftest_perfCtrl_dump,
  input  [63:0] difftest_logCtrl_begin,
  input  [63:0] difftest_logCtrl_end,
  input  [63:0] difftest_logCtrl_level,
  output        difftest_uart_out_valid,
  output [7:0]  difftest_uart_out_ch,
  output        difftest_uart_in_valid,
  input  [7:0]  difftest_uart_in_ch
);

  wire         _jtag_jtag_TCK;
  wire         _jtag_jtag_TMS;
  wire         _jtag_jtag_TDI;
  wire         _memory_io_axi4_0_aw_ready;
  wire         _memory_io_axi4_0_w_ready;
  wire         _memory_io_axi4_0_b_valid;
  wire [13:0]  _memory_io_axi4_0_b_bits_id;
  wire [1:0]   _memory_io_axi4_0_b_bits_resp;
  wire         _memory_io_axi4_0_ar_ready;
  wire         _memory_io_axi4_0_r_valid;
  wire [13:0]  _memory_io_axi4_0_r_bits_id;
  wire [255:0] _memory_io_axi4_0_r_bits_data;
  wire [1:0]   _memory_io_axi4_0_r_bits_resp;
  wire         _memory_io_axi4_0_r_bits_last;
  wire         _l_simMMIO_io_axi4_0_aw_ready;
  wire         _l_simMMIO_io_axi4_0_w_ready;
  wire         _l_simMMIO_io_axi4_0_b_valid;
  wire [1:0]   _l_simMMIO_io_axi4_0_b_bits_id;
  wire [1:0]   _l_simMMIO_io_axi4_0_b_bits_resp;
  wire         _l_simMMIO_io_axi4_0_ar_ready;
  wire         _l_simMMIO_io_axi4_0_r_valid;
  wire [1:0]   _l_simMMIO_io_axi4_0_r_bits_id;
  wire [63:0]  _l_simMMIO_io_axi4_0_r_bits_data;
  wire [1:0]   _l_simMMIO_io_axi4_0_r_bits_resp;
  wire         _l_simMMIO_io_axi4_0_r_bits_last;
  wire [63:0]  _l_simMMIO_io_interrupt_intrVec;
  wire         _l_soc_peripheral_awvalid;
  wire [1:0]   _l_soc_peripheral_awid;
  wire [30:0]  _l_soc_peripheral_awaddr;
  wire [7:0]   _l_soc_peripheral_awlen;
  wire [2:0]   _l_soc_peripheral_awsize;
  wire [1:0]   _l_soc_peripheral_awburst;
  wire         _l_soc_peripheral_awlock;
  wire [3:0]   _l_soc_peripheral_awcache;
  wire [2:0]   _l_soc_peripheral_awprot;
  wire [3:0]   _l_soc_peripheral_awqos;
  wire         _l_soc_peripheral_wvalid;
  wire [63:0]  _l_soc_peripheral_wdata;
  wire [7:0]   _l_soc_peripheral_wstrb;
  wire         _l_soc_peripheral_wlast;
  wire         _l_soc_peripheral_bready;
  wire         _l_soc_peripheral_arvalid;
  wire [1:0]   _l_soc_peripheral_arid;
  wire [30:0]  _l_soc_peripheral_araddr;
  wire [7:0]   _l_soc_peripheral_arlen;
  wire [2:0]   _l_soc_peripheral_arsize;
  wire [1:0]   _l_soc_peripheral_arburst;
  wire         _l_soc_peripheral_arlock;
  wire [3:0]   _l_soc_peripheral_arcache;
  wire [2:0]   _l_soc_peripheral_arprot;
  wire [3:0]   _l_soc_peripheral_arqos;
  wire         _l_soc_peripheral_rready;
  wire         _l_soc_memory_awvalid;
  wire [13:0]  _l_soc_memory_awid;
  wire [47:0]  _l_soc_memory_awaddr;
  wire [7:0]   _l_soc_memory_awlen;
  wire [2:0]   _l_soc_memory_awsize;
  wire [1:0]   _l_soc_memory_awburst;
  wire         _l_soc_memory_awlock;
  wire [3:0]   _l_soc_memory_awcache;
  wire [2:0]   _l_soc_memory_awprot;
  wire [3:0]   _l_soc_memory_awqos;
  wire         _l_soc_memory_wvalid;
  wire [255:0] _l_soc_memory_wdata;
  wire [31:0]  _l_soc_memory_wstrb;
  wire         _l_soc_memory_wlast;
  wire         _l_soc_memory_bready;
  wire         _l_soc_memory_arvalid;
  wire [13:0]  _l_soc_memory_arid;
  wire [47:0]  _l_soc_memory_araddr;
  wire [7:0]   _l_soc_memory_arlen;
  wire [2:0]   _l_soc_memory_arsize;
  wire [1:0]   _l_soc_memory_arburst;
  wire         _l_soc_memory_arlock;
  wire [3:0]   _l_soc_memory_arcache;
  wire [2:0]   _l_soc_memory_arprot;
  wire [3:0]   _l_soc_memory_arqos;
  wire         _l_soc_memory_rready;
  wire         _l_soc_io_systemjtag_jtag_TDO_data;
  wire         _l_soc_io_systemjtag_jtag_TDO_driven;
  wire         _l_soc_io_debug_reset;
  reg  [5:0]   rtcCounter;
  reg          rtcClock;
  reg  [63:0]  difftest_timer;
  wire         difftest_log_enable =
    difftest_timer >= difftest_logCtrl_begin & difftest_timer < difftest_logCtrl_end;
  always @(posedge clock) begin
    if (reset) begin
      rtcCounter <= 6'h0;
      rtcClock <= 1'h0;
      difftest_timer <= 64'h0;
    end
    else begin
      if (rtcCounter == 6'h31)
        rtcCounter <= 6'h0;
      else
        rtcCounter <= 6'(rtcCounter + 6'h1);
      rtcClock <= rtcCounter == 6'h0 ^ rtcClock;
      difftest_timer <= 64'(difftest_timer + 64'h1);
    end
  end // always @(posedge)
  `ifdef ENABLE_INITIAL_REG_
    `ifdef FIRRTL_BEFORE_INITIAL
      `FIRRTL_BEFORE_INITIAL
    `endif // FIRRTL_BEFORE_INITIAL
    logic [31:0] _RANDOM[0:2];
    initial begin
      `ifdef INIT_RANDOM_PROLOG_
        `INIT_RANDOM_PROLOG_
      `endif // INIT_RANDOM_PROLOG_
      `ifdef RANDOMIZE_REG_INIT
        for (logic [1:0] i = 2'h0; i < 2'h3; i += 2'h1) begin
          _RANDOM[i] = `RANDOM;
        end
        rtcCounter = _RANDOM[2'h0][5:0];
        rtcClock = _RANDOM[2'h0][6];
        difftest_timer = {_RANDOM[2'h0][31:7], _RANDOM[2'h1], _RANDOM[2'h2][6:0]};
      `endif // RANDOMIZE_REG_INIT
    end // initial
    `ifdef FIRRTL_AFTER_INITIAL
      `FIRRTL_AFTER_INITIAL
    `endif // FIRRTL_AFTER_INITIAL
  `endif // ENABLE_INITIAL_REG_
  XSTop l_soc (
    .nmi_0_0                                     (1'h0),
    .nmi_0_1                                     (1'h0),
    .dma_awready                                 (/* unused */),
    .dma_awvalid                                 (1'h0),
    .dma_awid                                    (14'h0),
    .dma_awaddr                                  (48'h0),
    .dma_awlen                                   (8'h0),
    .dma_awsize                                  (3'h0),
    .dma_awburst                                 (2'h0),
    .dma_awlock                                  (1'h0),
    .dma_awcache                                 (4'h0),
    .dma_awprot                                  (3'h0),
    .dma_awqos                                   (4'h0),
    .dma_wready                                  (/* unused */),
    .dma_wvalid                                  (1'h0),
    .dma_wdata                                   (256'h0),
    .dma_wstrb                                   (32'h0),
    .dma_wlast                                   (1'h0),
    .dma_bready                                  (1'h0),
    .dma_bvalid                                  (/* unused */),
    .dma_bid                                     (/* unused */),
    .dma_bresp                                   (/* unused */),
    .dma_arready                                 (/* unused */),
    .dma_arvalid                                 (1'h0),
    .dma_arid                                    (14'h0),
    .dma_araddr                                  (48'h0),
    .dma_arlen                                   (8'h0),
    .dma_arsize                                  (3'h0),
    .dma_arburst                                 (2'h0),
    .dma_arlock                                  (1'h0),
    .dma_arcache                                 (4'h0),
    .dma_arprot                                  (3'h0),
    .dma_arqos                                   (4'h0),
    .dma_rready                                  (1'h0),
    .dma_rvalid                                  (/* unused */),
    .dma_rid                                     (/* unused */),
    .dma_rdata                                   (/* unused */),
    .dma_rresp                                   (/* unused */),
    .dma_rlast                                   (/* unused */),
    .peripheral_awready                          (_l_simMMIO_io_axi4_0_aw_ready),
    .peripheral_awvalid                          (_l_soc_peripheral_awvalid),
    .peripheral_awid                             (_l_soc_peripheral_awid),
    .peripheral_awaddr                           (_l_soc_peripheral_awaddr),
    .peripheral_awlen                            (_l_soc_peripheral_awlen),
    .peripheral_awsize                           (_l_soc_peripheral_awsize),
    .peripheral_awburst                          (_l_soc_peripheral_awburst),
    .peripheral_awlock                           (_l_soc_peripheral_awlock),
    .peripheral_awcache                          (_l_soc_peripheral_awcache),
    .peripheral_awprot                           (_l_soc_peripheral_awprot),
    .peripheral_awqos                            (_l_soc_peripheral_awqos),
    .peripheral_wready                           (_l_simMMIO_io_axi4_0_w_ready),
    .peripheral_wvalid                           (_l_soc_peripheral_wvalid),
    .peripheral_wdata                            (_l_soc_peripheral_wdata),
    .peripheral_wstrb                            (_l_soc_peripheral_wstrb),
    .peripheral_wlast                            (_l_soc_peripheral_wlast),
    .peripheral_bready                           (_l_soc_peripheral_bready),
    .peripheral_bvalid                           (_l_simMMIO_io_axi4_0_b_valid),
    .peripheral_bid                              (_l_simMMIO_io_axi4_0_b_bits_id),
    .peripheral_bresp                            (_l_simMMIO_io_axi4_0_b_bits_resp),
    .peripheral_arready                          (_l_simMMIO_io_axi4_0_ar_ready),
    .peripheral_arvalid                          (_l_soc_peripheral_arvalid),
    .peripheral_arid                             (_l_soc_peripheral_arid),
    .peripheral_araddr                           (_l_soc_peripheral_araddr),
    .peripheral_arlen                            (_l_soc_peripheral_arlen),
    .peripheral_arsize                           (_l_soc_peripheral_arsize),
    .peripheral_arburst                          (_l_soc_peripheral_arburst),
    .peripheral_arlock                           (_l_soc_peripheral_arlock),
    .peripheral_arcache                          (_l_soc_peripheral_arcache),
    .peripheral_arprot                           (_l_soc_peripheral_arprot),
    .peripheral_arqos                            (_l_soc_peripheral_arqos),
    .peripheral_rready                           (_l_soc_peripheral_rready),
    .peripheral_rvalid                           (_l_simMMIO_io_axi4_0_r_valid),
    .peripheral_rid                              (_l_simMMIO_io_axi4_0_r_bits_id),
    .peripheral_rdata                            (_l_simMMIO_io_axi4_0_r_bits_data),
    .peripheral_rresp                            (_l_simMMIO_io_axi4_0_r_bits_resp),
    .peripheral_rlast                            (_l_simMMIO_io_axi4_0_r_bits_last),
    .memory_awready                              (_memory_io_axi4_0_aw_ready),
    .memory_awvalid                              (_l_soc_memory_awvalid),
    .memory_awid                                 (_l_soc_memory_awid),
    .memory_awaddr                               (_l_soc_memory_awaddr),
    .memory_awlen                                (_l_soc_memory_awlen),
    .memory_awsize                               (_l_soc_memory_awsize),
    .memory_awburst                              (_l_soc_memory_awburst),
    .memory_awlock                               (_l_soc_memory_awlock),
    .memory_awcache                              (_l_soc_memory_awcache),
    .memory_awprot                               (_l_soc_memory_awprot),
    .memory_awqos                                (_l_soc_memory_awqos),
    .memory_wready                               (_memory_io_axi4_0_w_ready),
    .memory_wvalid                               (_l_soc_memory_wvalid),
    .memory_wdata                                (_l_soc_memory_wdata),
    .memory_wstrb                                (_l_soc_memory_wstrb),
    .memory_wlast                                (_l_soc_memory_wlast),
    .memory_bready                               (_l_soc_memory_bready),
    .memory_bvalid                               (_memory_io_axi4_0_b_valid),
    .memory_bid                                  (_memory_io_axi4_0_b_bits_id),
    .memory_bresp                                (_memory_io_axi4_0_b_bits_resp),
    .memory_arready                              (_memory_io_axi4_0_ar_ready),
    .memory_arvalid                              (_l_soc_memory_arvalid),
    .memory_arid                                 (_l_soc_memory_arid),
    .memory_araddr                               (_l_soc_memory_araddr),
    .memory_arlen                                (_l_soc_memory_arlen),
    .memory_arsize                               (_l_soc_memory_arsize),
    .memory_arburst                              (_l_soc_memory_arburst),
    .memory_arlock                               (_l_soc_memory_arlock),
    .memory_arcache                              (_l_soc_memory_arcache),
    .memory_arprot                               (_l_soc_memory_arprot),
    .memory_arqos                                (_l_soc_memory_arqos),
    .memory_rready                               (_l_soc_memory_rready),
    .memory_rvalid                               (_memory_io_axi4_0_r_valid),
    .memory_rid                                  (_memory_io_axi4_0_r_bits_id),
    .memory_rdata                                (_memory_io_axi4_0_r_bits_data),
    .memory_rresp                                (_memory_io_axi4_0_r_bits_resp),
    .memory_rlast                                (_memory_io_axi4_0_r_bits_last),
    .io_clock                                    (clock),
    .io_reset                                    (reset | _l_soc_io_debug_reset),
    .io_sram_config                              (16'h0),
    .io_extIntrs                                 (_l_simMMIO_io_interrupt_intrVec),
    .io_pll0_lock                                (1'h1),
    .io_pll0_ctrl_0                              (/* unused */),
    .io_pll0_ctrl_1                              (/* unused */),
    .io_pll0_ctrl_2                              (/* unused */),
    .io_pll0_ctrl_3                              (/* unused */),
    .io_pll0_ctrl_4                              (/* unused */),
    .io_pll0_ctrl_5                              (/* unused */),
    .io_systemjtag_jtag_TCK                      (_jtag_jtag_TCK),
    .io_systemjtag_jtag_TMS                      (_jtag_jtag_TMS),
    .io_systemjtag_jtag_TDI                      (_jtag_jtag_TDI),
    .io_systemjtag_jtag_TDO_data                 (_l_soc_io_systemjtag_jtag_TDO_data),
    .io_systemjtag_jtag_TDO_driven               (_l_soc_io_systemjtag_jtag_TDO_driven),
    .io_systemjtag_reset                         (reset),
    .io_systemjtag_mfr_id                        (11'h0),
    .io_systemjtag_part_number                   (16'h0),
    .io_systemjtag_version                       (4'h0),
    .io_debug_reset                              (_l_soc_io_debug_reset),
    .io_rtc_clock                                (rtcClock),
    .io_cacheable_check_req_0_valid              (1'h0),
    .io_cacheable_check_req_0_bits_addr          (48'h0),
    .io_cacheable_check_req_0_bits_size          (2'h0),
    .io_cacheable_check_req_0_bits_cmd           (3'h0),
    .io_cacheable_check_req_1_valid              (1'h0),
    .io_cacheable_check_req_1_bits_addr          (48'h0),
    .io_cacheable_check_req_1_bits_size          (2'h0),
    .io_cacheable_check_req_1_bits_cmd           (3'h0),
    .io_cacheable_check_resp_0_ld                (/* unused */),
    .io_cacheable_check_resp_0_st                (/* unused */),
    .io_cacheable_check_resp_0_instr             (/* unused */),
    .io_cacheable_check_resp_0_mmio              (/* unused */),
    .io_cacheable_check_resp_0_atomic            (/* unused */),
    .io_cacheable_check_resp_1_ld                (/* unused */),
    .io_cacheable_check_resp_1_st                (/* unused */),
    .io_cacheable_check_resp_1_instr             (/* unused */),
    .io_cacheable_check_resp_1_mmio              (/* unused */),
    .io_cacheable_check_resp_1_atomic            (/* unused */),
    .io_riscv_halt_0                             (/* unused */),
    .io_riscv_critical_error_0                   (/* unused */),
    .io_riscv_rst_vec_0                          (48'h10000000),
    .io_traceCoreInterface_0_fromEncoder_enable  (1'h0),
    .io_traceCoreInterface_0_fromEncoder_stall   (1'h0),
    .io_traceCoreInterface_0_toEncoder_cause     (/* unused */),
    .io_traceCoreInterface_0_toEncoder_tval      (/* unused */),
    .io_traceCoreInterface_0_toEncoder_priv      (/* unused */),
    .io_traceCoreInterface_0_toEncoder_iaddr     (/* unused */),
    .io_traceCoreInterface_0_toEncoder_itype     (/* unused */),
    .io_traceCoreInterface_0_toEncoder_iretire   (/* unused */),
    .io_traceCoreInterface_0_toEncoder_ilastsize (/* unused */)
  );
  SimMMIO l_simMMIO (
    .clock                   (clock),
    .reset                   (reset),
    .io_axi4_0_aw_ready      (_l_simMMIO_io_axi4_0_aw_ready),
    .io_axi4_0_aw_valid      (_l_soc_peripheral_awvalid),
    .io_axi4_0_aw_bits_id    (_l_soc_peripheral_awid),
    .io_axi4_0_aw_bits_addr  (_l_soc_peripheral_awaddr),
    .io_axi4_0_aw_bits_len   (_l_soc_peripheral_awlen),
    .io_axi4_0_aw_bits_size  (_l_soc_peripheral_awsize),
    .io_axi4_0_aw_bits_burst (_l_soc_peripheral_awburst),
    .io_axi4_0_aw_bits_lock  (_l_soc_peripheral_awlock),
    .io_axi4_0_aw_bits_cache (_l_soc_peripheral_awcache),
    .io_axi4_0_aw_bits_prot  (_l_soc_peripheral_awprot),
    .io_axi4_0_aw_bits_qos   (_l_soc_peripheral_awqos),
    .io_axi4_0_w_ready       (_l_simMMIO_io_axi4_0_w_ready),
    .io_axi4_0_w_valid       (_l_soc_peripheral_wvalid),
    .io_axi4_0_w_bits_data   (_l_soc_peripheral_wdata),
    .io_axi4_0_w_bits_strb   (_l_soc_peripheral_wstrb),
    .io_axi4_0_w_bits_last   (_l_soc_peripheral_wlast),
    .io_axi4_0_b_ready       (_l_soc_peripheral_bready),
    .io_axi4_0_b_valid       (_l_simMMIO_io_axi4_0_b_valid),
    .io_axi4_0_b_bits_id     (_l_simMMIO_io_axi4_0_b_bits_id),
    .io_axi4_0_b_bits_resp   (_l_simMMIO_io_axi4_0_b_bits_resp),
    .io_axi4_0_ar_ready      (_l_simMMIO_io_axi4_0_ar_ready),
    .io_axi4_0_ar_valid      (_l_soc_peripheral_arvalid),
    .io_axi4_0_ar_bits_id    (_l_soc_peripheral_arid),
    .io_axi4_0_ar_bits_addr  (_l_soc_peripheral_araddr),
    .io_axi4_0_ar_bits_len   (_l_soc_peripheral_arlen),
    .io_axi4_0_ar_bits_size  (_l_soc_peripheral_arsize),
    .io_axi4_0_ar_bits_burst (_l_soc_peripheral_arburst),
    .io_axi4_0_ar_bits_lock  (_l_soc_peripheral_arlock),
    .io_axi4_0_ar_bits_cache (_l_soc_peripheral_arcache),
    .io_axi4_0_ar_bits_prot  (_l_soc_peripheral_arprot),
    .io_axi4_0_ar_bits_qos   (_l_soc_peripheral_arqos),
    .io_axi4_0_r_ready       (_l_soc_peripheral_rready),
    .io_axi4_0_r_valid       (_l_simMMIO_io_axi4_0_r_valid),
    .io_axi4_0_r_bits_id     (_l_simMMIO_io_axi4_0_r_bits_id),
    .io_axi4_0_r_bits_data   (_l_simMMIO_io_axi4_0_r_bits_data),
    .io_axi4_0_r_bits_resp   (_l_simMMIO_io_axi4_0_r_bits_resp),
    .io_axi4_0_r_bits_last   (_l_simMMIO_io_axi4_0_r_bits_last),
    .io_uart_out_valid       (difftest_uart_out_valid),
    .io_uart_out_ch          (difftest_uart_out_ch),
    .io_uart_in_valid        (difftest_uart_in_valid),
    .io_uart_in_ch           (difftest_uart_in_ch),
    .io_interrupt_intrVec    (_l_simMMIO_io_interrupt_intrVec)
  );
  AXI4RAMWrapper memory (
    .clock                   (clock),
    .reset                   (reset),
    .io_axi4_0_aw_ready      (_memory_io_axi4_0_aw_ready),
    .io_axi4_0_aw_valid      (_l_soc_memory_awvalid),
    .io_axi4_0_aw_bits_id    (_l_soc_memory_awid),
    .io_axi4_0_aw_bits_addr  (_l_soc_memory_awaddr),
    .io_axi4_0_aw_bits_len   (_l_soc_memory_awlen),
    .io_axi4_0_aw_bits_size  (_l_soc_memory_awsize),
    .io_axi4_0_aw_bits_burst (_l_soc_memory_awburst),
    .io_axi4_0_aw_bits_lock  (_l_soc_memory_awlock),
    .io_axi4_0_aw_bits_cache (_l_soc_memory_awcache),
    .io_axi4_0_aw_bits_prot  (_l_soc_memory_awprot),
    .io_axi4_0_aw_bits_qos   (_l_soc_memory_awqos),
    .io_axi4_0_w_ready       (_memory_io_axi4_0_w_ready),
    .io_axi4_0_w_valid       (_l_soc_memory_wvalid),
    .io_axi4_0_w_bits_data   (_l_soc_memory_wdata),
    .io_axi4_0_w_bits_strb   (_l_soc_memory_wstrb),
    .io_axi4_0_w_bits_last   (_l_soc_memory_wlast),
    .io_axi4_0_b_ready       (_l_soc_memory_bready),
    .io_axi4_0_b_valid       (_memory_io_axi4_0_b_valid),
    .io_axi4_0_b_bits_id     (_memory_io_axi4_0_b_bits_id),
    .io_axi4_0_b_bits_resp   (_memory_io_axi4_0_b_bits_resp),
    .io_axi4_0_ar_ready      (_memory_io_axi4_0_ar_ready),
    .io_axi4_0_ar_valid      (_l_soc_memory_arvalid),
    .io_axi4_0_ar_bits_id    (_l_soc_memory_arid),
    .io_axi4_0_ar_bits_addr  (_l_soc_memory_araddr),
    .io_axi4_0_ar_bits_len   (_l_soc_memory_arlen),
    .io_axi4_0_ar_bits_size  (_l_soc_memory_arsize),
    .io_axi4_0_ar_bits_burst (_l_soc_memory_arburst),
    .io_axi4_0_ar_bits_lock  (_l_soc_memory_arlock),
    .io_axi4_0_ar_bits_cache (_l_soc_memory_arcache),
    .io_axi4_0_ar_bits_prot  (_l_soc_memory_arprot),
    .io_axi4_0_ar_bits_qos   (_l_soc_memory_arqos),
    .io_axi4_0_r_ready       (_l_soc_memory_rready),
    .io_axi4_0_r_valid       (_memory_io_axi4_0_r_valid),
    .io_axi4_0_r_bits_id     (_memory_io_axi4_0_r_bits_id),
    .io_axi4_0_r_bits_data   (_memory_io_axi4_0_r_bits_data),
    .io_axi4_0_r_bits_resp   (_memory_io_axi4_0_r_bits_resp),
    .io_axi4_0_r_bits_last   (_memory_io_axi4_0_r_bits_last)
  );
  SimJTAG #(
    .TICK_DELAY(3)
  ) jtag (
    .clock           (clock),
    .reset           (reset),
    .jtag_TRSTn      (/* unused */),
    .jtag_TCK        (_jtag_jtag_TCK),
    .jtag_TMS        (_jtag_jtag_TMS),
    .jtag_TDI        (_jtag_jtag_TDI),
    .jtag_TDO_data   (_l_soc_io_systemjtag_jtag_TDO_data),
    .jtag_TDO_driven (_l_soc_io_systemjtag_jtag_TDO_driven),
    .enable          (1'h1),
    .init_done       (~reset),
    .exit            (/* unused */)
  );
  assign difftest_exit = 64'h0;
  assign difftest_step = 64'h1;
endmodule

