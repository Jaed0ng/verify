module tb_top;
  `include "xs_tests.svh"

  // 实例化接口
  xs_top_if vif();

  // 实例化DUT
  XSTop dut (
    .nmi_0_0                     (vif.nmi_0_0),
    .nmi_0_1                     (vif.nmi_0_1),
    .dma_awready                 (vif.dma_awready),
    .dma_awvalid                 (vif.dma_awvalid),
    .dma_awid                    (vif.dma_awid),
    .dma_awaddr                  (vif.dma_awaddr),
    .dma_awlen                   (vif.dma_awlen),
    .dma_awsize                  (vif.dma_awsize),
    .dma_awburst                 (vif.dma_awburst),
    .dma_awlock                  (vif.dma_awlock),
    .dma_awcache                 (vif.dma_awcache),
    .dma_awprot                  (vif.dma_awprot),
    .dma_awqos                   (vif.dma_awqos),
    .dma_wready                  (vif.dma_wready),
    .dma_wvalid                  (vif.dma_wvalid),
    .dma_wdata                   (vif.dma_wdata),
    .dma_wstrb                   (vif.dma_wstrb),
    .dma_wlast                   (vif.dma_wlast),
    .dma_bready                  (vif.dma_bready),
    .dma_bvalid                  (vif.dma_bvalid),
    .dma_bid                     (vif.dma_bid),
    .dma_bresp                   (vif.dma_bresp),
    .dma_arready                 (vif.dma_arready),
    .dma_arvalid                 (vif.dma_arvalid),
    .dma_arid                    (vif.dma_arid),
    .dma_araddr                  (vif.dma_araddr),
    .dma_arlen                   (vif.dma_arlen),
    .dma_arsize                  (vif.dma_arsize),
    .dma_arburst                 (vif.dma_arburst),
    .dma_arlock                  (vif.dma_arlock),
    .dma_arcache                 (vif.dma_arcache),
    .dma_arprot                  (vif.dma_arprot),
    .dma_arqos                   (vif.dma_arqos),
    .dma_rready                  (vif.dma_rready),
    .dma_rvalid                  (vif.dma_rvalid),
    .dma_rid                     (vif.dma_rid),
    .dma_rdata                   (vif.dma_rdata),
    .dma_rresp                   (vif.dma_rresp),
    .dma_rlast                   (vif.dma_rlast),
    .peripheral_awready          (vif.peripheral_awready),
    .peripheral_awvalid          (vif.peripheral_awvalid),
    .peripheral_awid             (vif.peripheral_awid),
    .peripheral_awaddr           (vif.peripheral_awaddr),
    .peripheral_awlen            (vif.peripheral_awlen),
    .peripheral_awsize           (vif.peripheral_awsize),
    .peripheral_awburst          (vif.peripheral_awburst),
    .peripheral_awlock           (vif.peripheral_awlock),
    .peripheral_awcache          (vif.peripheral_awcache),
    .peripheral_awprot           (vif.peripheral_awprot),
    .peripheral_awqos            (vif.peripheral_awqos),
    .peripheral_wready           (vif.peripheral_wready),
    .peripheral_wvalid           (vif.peripheral_wvalid),
    .peripheral_wdata            (vif.peripheral_wdata),
    .peripheral_wstrb            (vif.peripheral_wstrb),
    .peripheral_wlast            (vif.peripheral_wlast),
    .peripheral_bready           (vif.peripheral_bready),
    .peripheral_bvalid           (vif.peripheral_bvalid),
    .peripheral_bid              (vif.peripheral_bid),
    .peripheral_bresp            (vif.peripheral_bresp),
    .peripheral_arready          (vif.peripheral_arready),
    .peripheral_arvalid          (vif.peripheral_arvalid),
    .peripheral_arid             (vif.peripheral_arid),
    .peripheral_araddr           (vif.peripheral_araddr),
    .peripheral_arlen            (vif.peripheral_arlen),
    .peripheral_arsize           (vif.peripheral_arsize),
    .peripheral_arburst          (vif.peripheral_arburst),
    .peripheral_arlock           (vif.peripheral_arlock),
    .peripheral_arcache          (vif.peripheral_arcache),
    .peripheral_arprot           (vif.peripheral_arprot),
    .peripheral_arqos            (vif.peripheral_arqos),
    .peripheral_rready           (vif.peripheral_rready),
    .peripheral_rvalid           (vif.peripheral_rvalid),
    .peripheral_rid              (vif.peripheral_rid),
    .peripheral_rdata            (vif.peripheral_rdata),
    .peripheral_rresp            (vif.peripheral_rresp),
    .peripheral_rlast            (vif.peripheral_rlast),
    .memory_awready              (vif.memory_awready),
    .memory_awvalid              (vif.memory_awvalid),
    .memory_awid                 (vif.memory_awid),
    .memory_awaddr               (vif.memory_awaddr),
    .memory_awlen                (vif.memory_awlen),
    .memory_awsize               (vif.memory_awsize),
    .memory_awburst              (vif.memory_awburst),
    .memory_awlock               (vif.memory_awlock),
    .memory_awcache              (vif.memory_awcache),
    .memory_awprot               (vif.memory_awprot),
    .memory_awqos                (vif.memory_awqos),
    .memory_wready               (vif.memory_wready),
    .memory_wvalid               (vif.memory_wvalid),
    .memory_wdata                (vif.memory_wdata),
    .memory_wstrb                (vif.memory_wstrb),
    .memory_wlast                (vif.memory_wlast),
    .memory_bready               (vif.memory_bready),
    .memory_bvalid               (vif.memory_bvalid),
    .memory_bid                  (vif.memory_bid),
    .memory_bresp                (vif.memory_bresp),
    .memory_arready              (vif.memory_arready),
    .memory_arvalid              (vif.memory_arvalid),
    .memory_arid                 (vif.memory_arid),
    .memory_araddr               (vif.memory_araddr),
    .memory_arlen                (vif.memory_arlen),
    .memory_arsize               (vif.memory_arsize),
    .memory_arburst              (vif.memory_arburst),
    .memory_arlock               (vif.memory_arlock),
    .memory_arcache              (vif.memory_arcache),
    .memory_arprot               (vif.memory_arprot),
    .memory_arqos                (vif.memory_arqos),
    .memory_rready               (vif.memory_rready),
    .memory_rvalid               (vif.memory_rvalid),
    .memory_rid                  (vif.memory_rid),
    .memory_rdata                (vif.memory_rdata),
    .memory_rresp                (vif.memory_rresp),
    .memory_rlast                (vif.memory_rlast),
    .io_clock                    (vif.io_clock),
    .io_reset                    (vif.io_reset),
    .io_sram_config              (vif.io_sram_config),
    .io_extIntrs                 (vif.io_extIntrs),
    .io_pll0_lock                (vif.io_pll0_lock),
    .io_pll0_ctrl_0              (vif.io_pll0_ctrl_0),
    .io_pll0_ctrl_1              (vif.io_pll0_ctrl_1),
    .io_pll0_ctrl_2              (vif.io_pll0_ctrl_2),
    .io_pll0_ctrl_3              (vif.io_pll0_ctrl_3),
    .io_pll0_ctrl_4              (vif.io_pll0_ctrl_4),
    .io_pll0_ctrl_5              (vif.io_pll0_ctrl_5),
    .io_systemjtag_jtag_TCK      (vif.io_systemjtag_jtag_TCK),
    .io_systemjtag_jtag_TMS      (vif.io_systemjtag_jtag_TMS),
    .io_systemjtag_jtag_TDI      (vif.io_systemjtag_jtag_TDI),
    .io_systemjtag_jtag_TDO_data (vif.io_systemjtag_jtag_TDO_data),
    .io_systemjtag_jtag_TDO_driven (vif.io_systemjtag_jtag_TDO_driven),
    .io_systemjtag_reset         (vif.io_systemjtag_reset),
    .io_systemjtag_mfr_id        (vif.io_systemjtag_mfr_id),
    .io_systemjtag_part_number   (vif.io_systemjtag_part_number),
    .io_systemjtag_version       (vif.io_systemjtag_version),
    .io_debug_reset              (vif.io_debug_reset),
    .io_rtc_clock                (vif.io_rtc_clock),
    .io_cacheable_check_req_0_valid (1'b0),
    .io_cacheable_check_req_0_bits_addr (48'h0),
    .io_cacheable_check_req_0_bits_size (2'h0),
    .io_cacheable_check_req_0_bits_cmd (3'h0),
    .io_cacheable_check_req_1_valid (1'b0),
    .io_cacheable_check_req_1_bits_addr (48'h0),
    .io_cacheable_check_req_1_bits_size (2'h0),
    .io_cacheable_check_req_1_bits_cmd (3'h0),
    .io_riscv_halt_0             (vif.io_riscv_halt_0),
    .io_riscv_critical_error_0   (vif.io_riscv_critical_error_0),
    .io_riscv_rst_vec_0          (vif.io_riscv_rst_vec_0),
    .io_traceCoreInterface_0_fromEncoder_enable (1'b0),
    .io_traceCoreInterface_0_fromEncoder_stall (1'b0)
  );

  // 配置UVM并启动仿真
  initial begin
    // 注册接口到UVM配置数据库
    uvm_config_db#(virtual xs_top_if)::set(null, "*", "vif", vif);
    // 启动UVM仿真
    run_test("");
  end

  // 生成波形文件
  initial begin         
    $fsdbDumpfile("tb_top.fsdb");
    $fsdbDumpvars(0,tb_top); 
  end

endmodule

